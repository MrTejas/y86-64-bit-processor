`include "ANDx64.v"
module ANDx64_test();

reg signed [63:0] a;
reg signed [63:0] b;

wire signed [63:0] ans;

ANDx64 AT23(a,b,ans);

initial
    begin
        $dumpfile("ANDx64_test.vcd");
        $dumpvars(0, ANDx64_test);
        a = 64'b0;
        b = 64'b0;
        
        $monitor("time: %0d\n a  : %b\t%d\n b  : %b\t%d\n ans: %b\t%d\n", $time, a,a,b,b,ans,ans);

        // #5 a = 64'd2811; b= 64'd1012;
        // #5 a = -64'd1243; b= 64'd1234;
        // #5 a = -64'd7478; b=-64'd46474;
        // #5 a = 64'd1092835; b = -64'd1020;
        // #5 a = 64'd7890678653; b = 64'd4238598110567;
        // #5 a = 64'b0111111111111111111111111111111111111111111111111111111111111111; b = 64'd1;
        // #5 a = -64'd9223372036854770000; b=-64'd6000;
        // #5 a = 64'd4238; b=-64'd4238;
        // #5 a = -64'd4238598110567; b = -64'd4238598110567;

        // edge cases
        
        #5 a = -64'd9223372036854775808; b = -64'd9223372036854775808;
        #5 a = 64'd9223372036854775807; b = 64'd9223372036854775807;
        #5 a = 64'd9223372036854775807; b = -64'd9223372036854775808;
        #5 a = -64'd1; b = -64'd9223372036854775808;
    end
endmodule