`timescale 10ps/1ps
`include "SUBx1.v"
`include "SUBx64.v"

module tb_SUBx64();

reg signed [63:0] a;
reg signed [63:0] b;

wire signed [63:0] diff;
wire OF;

SUBx64 AT22(a,b,diff,OF);

initial
    begin
        $dumpfile("tb_SUBx64.vcd");
        $dumpvars(0, tb_SUBx64);
        a = 64'b0;
        b = 64'b0;
        
        $monitor("time: %0d\n a  : %b\t%d\n b  : %b\t%d\n a-b: %b\t%d\n overflow=%b\n ", $time, a,a,b,b,diff,diff, OF);

        // #5 a = 64'd2811; b= 64'd1012;
        // #5 a = -64'd1243; b= 64'd1234;
        // #5 a = -64'd7478; b=-64'd46474;
        // #5 a = 64'd1092835; b = -64'd1020;
        // #5 a = 64'd7890678653; b = 64'd4238598110567;
        // #5 a = 64'b0111111111111111111111111111111111111111111111111111111111111111; b = 64'd1;
        // #5 a = -64'd9223372036854770000; b=-64'd6000;
        // #5 a = 64'd4238; b=-64'd4238;
        // #5 a = -64'd4238598110567; b = -64'd4238598110567;

        // // edge cases
        #10
        a = 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;
        b = 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;

        #10
        a = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
        b = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

        #10
        a = 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;
        b = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

        #10
        a = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
        b = 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;
        
    end
endmodule

// iverilog -o tb_SUBx64 tb_SUBx64.v
// vvp tb_SUBx64